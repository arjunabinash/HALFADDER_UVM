interface half_adder_if(input logic clk); 
  
  logic in_a;
  logic in_b;
  logic ena;
  logic sum;
  logic carry;
  
endinterface: half_adder_if